`timescale 1ns / 1ps

// Main algorithm to carry out decryption
// Module written and tested by C. Baldwin
module invMainAES(
    clk,
    aes_input,
    aes_key,
    aes_output      
    );
    
    // Declare inputs and outputs
    input clk;
    input [127:0] aes_input;
    input [127:0] aes_key;
    output [127:0] aes_output;
    
    // Declare other variables - these are the keys generated by the keyExpansion module and the outputs from each round
    wire [127:0] r0_key, r1_key, r2_key, r3_key, r4_key, r5_key, r6_key, r7_key, r8_key, r9_key, r10_key;
    wire [127:0] r0_output,  r1_output,  r2_output,  r3_output,  r4_output,  r5_output,  r6_output,  r7_output,  r8_output,  r9_output,  r10_output;
    
    // Generate 10 keys (key0 is the same as the initial cipher key)
    keyExpansion keys(clk, aes_key, r0_key, r1_key, r2_key, r3_key, r4_key, r5_key, r6_key, r7_key, r8_key, r9_key, r10_key);
    
    // Round 0 - simple XOR with initial cipher
    assign r0_output = aes_input^r10_key;
    
    // doRound function that carries out the operations for each round, passing the output to the next one
    doInvRound round1(clk, r0_output, r9_key, r1_output);
    doInvRound round2(clk, r1_output, r8_key, r2_output);
    doInvRound round3(clk, r2_output, r7_key, r3_output);
    doInvRound round4(clk, r3_output, r6_key, r4_output);
    doInvRound round5(clk, r4_output, r5_key, r5_output);
    doInvRound round6(clk, r5_output, r4_key, r6_output);
    doInvRound round7(clk, r6_output, r3_key, r7_output);
    doInvRound round8(clk, r7_output, r2_key, r8_output);
    doInvRound round9(clk, r8_output, r1_key, r9_output);
    // Final round - skips mix columns
    lastInvRound round10(clk, r9_output, r0_key, r10_output);
    
    // assign the output
    assign aes_output = r10_output;
    
endmodule
